ARCHITECTURE rtl OF vAdd IS
BEGIN
  sum <= sine +offset;
END rtl;
