ARCHITECTURE comb OF opConcatenate IS
BEGIN

  concatOut <= sine & concatIn;

END ARCHITECTURE comb;

