ARCHITECTURE comb OF opAdd IS
BEGIN

  sum <= sine + offset;

END ARCHITECTURE comb;

