ARCHITECTURE rtl OF vMultiply IS
BEGIN
  product <=sine * gain;
END rtl;
