ARCHITECTURE comb OF opMultiply IS
BEGIN

  product <= sine * gain;

END ARCHITECTURE comb;

