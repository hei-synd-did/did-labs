ARCHITECTURE studentVersion OF cordicStepAngles IS

BEGIN

  stepAngle0 <= "001000000000";
  stepAngle1 <= x"013";

END ARCHITECTURE studentVersion;
