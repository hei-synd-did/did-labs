ARCHITECTURE comb OF opInvert IS
BEGIN

  inverted <= not sine;

END ARCHITECTURE comb;

