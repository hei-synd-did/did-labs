ARCHITECTURE RTL OF vInvert IS
BEGIN
  inverted <= not sine;
END RTL;
