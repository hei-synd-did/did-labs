ARCHITECTURE rtl OF vConcatenate IS
BEGIN
  concatOut <= sine & concatIn;
END rtl;
